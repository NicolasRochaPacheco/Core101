


module DATA_MEM #(
  parameter XLEN = 32
)(
  input data_mem_valid_in,
  input data_mem_write_in,
  input [XLEN-1:0] data_mem_addr_in,
  input [XLEN-1:0] data_mem_data_in,
  output [XLEN-1:0] data_mem_data_out,
  output data_mem_ready_out
);




endmodule
