// Instruction memory module definition
// Copyright (C) 2019 Nicolas Rocha Pacheco
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <https://www.gnu.org/licenses/>.

module INS_MEM #(
  parameter XLEN = 32
)(
  input ins_mem_valid_in,
  input [XLEN-1:0] ins_mem_addr_in,
  output reg ins_mem_ready_out,
  output reg [XLEN-1:0] ins_mem_data_out
);

// Sets memory addressing width
parameter MEM_ADDR = 10;

// Parameter to set memory size
parameter MEM_SIZE = 2 ** MEM_ADDR;

// Defines memory
reg [7:0] ins_mem [0:MEM_SIZE-1];

initial
  $readmemh("./rtl/memory/ins_mem.hex", ins_mem);

always @ ( * ) begin
  if(ins_mem_valid_in == 1'b1) begin
    ins_mem_data_out = {
      ins_mem[ins_mem_addr_in[MEM_ADDR-1:0] + 3],
      ins_mem[ins_mem_addr_in[MEM_ADDR-1:0] + 2],
      ins_mem[ins_mem_addr_in[MEM_ADDR-1:0] + 1],
      ins_mem[ins_mem_addr_in[MEM_ADDR-1:0]]
    };
    ins_mem_ready_out = 1'b1;
  end
end

endmodule
