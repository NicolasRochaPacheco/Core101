module IMM_GEN(
  input   [31:0]  ins_input,
  output  [31:0]  imm_value_output
);


endmodule
