


module LSU_EXEC(
  input enable_in,
  input [31:0] a_data_in,
  input [31:0] b_data_in,

  output [31:0] res_data_out
);



endmodule
